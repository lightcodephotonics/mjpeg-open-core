// Copyright (c) 2018  LulinChen, All Rights Reserved
// AUTHOR : 	LulinChen
// AUTHOR'S EMAIL : lulinchen@aliyun.com 
// Release history
// VERSION Date AUTHOR DESCRIPTION
`include "jpeg_global.v"
module header_gen(
	input							clk,
	input 							rstn,	
	input 							header_go,	
	input							eoi,
	input     	[`W_PW:0]  			PicWidth_i,	
    input     	[`W_PH:0]  			PicHeight_i,	

	output reg						header_byte_f,
	output reg	[ 7:0]				header_byte,
	output reg						header_ready,
	output							frame_ready
	);
	//go	+|
	//max_f  					 +|
	//en	 |++++++++++++++++++++|
	//cnt	 |0..............MAX-1| MAX		
	reg					cnt_header_e;
	reg		[ 9:0]		cnt_header;
	wire				cnt_header_max_f = cnt_header == `HEADER_SIZE-1;
	always @(`CLK_RST_EDGE)
		if (`RST)					cnt_header_e <= 0;
		else if (header_go)			cnt_header_e <= 1;
		else if (cnt_header_max_f)	cnt_header_e <= 0;
	
	always @(`CLK_RST_EDGE)
		if (`RST)	cnt_header <= 0;
		else 		cnt_header <= cnt_header_e? cnt_header + 1 : 0;
	
	reg		[7:0]	cnt_header_e_d;
	always @(*)	cnt_header_e_d[0] = cnt_header_e;
	always @(`CLK_RST_EDGE)
		if (`RST)	cnt_header_e_d[7:1] <= 0;
		else 		cnt_header_e_d[7:1] <= cnt_header_e_d;
	reg		[7:0][9:0]	cnt_header_d;
	always @(*)	cnt_header_d[0] = cnt_header;
	always @(`CLK_RST_EDGE)
		if (`RST)	cnt_header_d[7:1] <= 0;
		else 		cnt_header_d[7:1] <= cnt_header_d;
	reg		[7:0]	cnt_header_max_f_d;
	always @(*)	cnt_header_max_f_d[0] = cnt_header_max_f;
	always @(`CLK_RST_EDGE)
		if (`RST)	cnt_header_max_f_d[7:1] <= 0;
		else 		cnt_header_max_f_d[7:1] <= cnt_header_max_f_d;	
		
	wire	[7:0]		q_rom_header;
	reg		[7:0]		q_rom_header_d1;
	always @(`CLK_RST_EDGE)
		if (`ZST)	q_rom_header_d1 <= 0;
		else 		q_rom_header_d1 <= q_rom_header;	
	
	// cnt  qa  qa_d1	header_byte_b1   header_byte
	reg				size_start;
	always @(`CLK_RST_EDGE)
		if (`RST)	size_start <= 0;
		else 		size_start <= cnt_header_d[1]== `ADDR_SIZE_Y_H;
	reg		[7:0]	size_start_d;
	always @(*)	size_start_d[0] = size_start;
	always @(`CLK_RST_EDGE)
		if (`RST)	size_start_d[7:1] <= 0;
		else 		size_start_d[7:1] <= size_start_d;	
	
	reg		[7:0]	header_byte_b1;
	always @(`CLK_RST_EDGE)
		if (`RST)					header_byte_b1 <= 0;
		else if (size_start)		header_byte_b1 <= PicHeight_i[`W_PH:8];
		else if (size_start_d[1])	header_byte_b1 <= PicHeight_i[7:0];
		else if (size_start_d[2])	header_byte_b1 <= PicWidth_i[`W_PW:8];
		else if (size_start_d[3])	header_byte_b1 <= PicWidth_i[7:0];
		else						header_byte_b1 <= q_rom_header_d1;
	
	rom_header rom_header(
		clk,
		cnt_header,
		q_rom_header
		);
	
	wire	[0:1][7:0]	EOI_bytes = 16'hFFD9;
	reg		eoi_e;
	always @(`CLK_RST_EDGE)
		if (`RST)	eoi_e <= 0;
		else 		eoi_e <= eoi;
	reg		[7:0]	eoi_e_d;
	always @(*)	eoi_e_d[0] = eoi_e;
	always @(`CLK_RST_EDGE)
		if (`RST)	eoi_e_d[7:1] <= 0;
		else 		eoi_e_d[7:1] <= eoi_e_d;
		
	assign	frame_ready = eoi_e_d[3];
	
	always @(`CLK_RST_EDGE)
		if (`RST)	header_byte_f <= 0;
		else 		header_byte_f <= cnt_header_e_d[3] | eoi_e | eoi_e_d[1];
	
	always @(`CLK_RST_EDGE)
		if (`RST)						header_byte <= 0;
		else if(cnt_header_e_d[3])		header_byte <= header_byte_b1;
		else if (eoi_e)					header_byte <= EOI_bytes[0];
		else if (eoi_e_d[1])			header_byte <= EOI_bytes[1];
	always @(`CLK_RST_EDGE)
		if (`RST)	header_ready <= 0;
		else 		header_ready <= cnt_header_max_f_d[3];
endmodule


module rom_header(
	input 				clk,
	input		[9:0]	addr,
	output reg	[7:0]	q
	);
	rom_header_qf09(clk,addr,q);
endmodule

module rom_header_qf02(
	input 				clk,
	input		[9:0]	addr,
	output reg	[7:0]	q
	);
	
	reg					[7:0]	rom [1023:0];
	always @(posedge clk) q <= rom[addr];
	initial begin
		rom[ 0    ] = 8'hFF;
		rom[ 1    ] = 8'hD8;
		rom[ 2    ] = 8'hFF;
		rom[ 3    ] = 8'hC0;
		rom[ 4    ] = 8'h00;
		rom[ 5    ] = 8'h11;
		rom[ 6    ] = 8'h08;
		rom[ 7    ] = 8'h01;
		rom[ 8    ] = 8'h20;
		rom[ 9    ] = 8'h01;
		rom[ 10   ] = 8'h60;
		rom[ 11   ] = 8'h03;
		rom[ 12   ] = 8'h01;
`ifdef YUV444_ONLY
		rom[ 13   ] = 8'h11;
`elsif YUV422_ONLY
		rom[ 13   ] = 8'h21;
`endif
		rom[ 14   ] = 8'h00;
		rom[ 15   ] = 8'h02;
		rom[ 16   ] = 8'h11;
		rom[ 17   ] = 8'h01;
		rom[ 18   ] = 8'h03;
		rom[ 19   ] = 8'h11;
		rom[ 20   ] = 8'h01;
		// quantization table index 0 header begins
		rom[ 21   ] = 8'hFF;
		rom[ 22   ] = 8'hDB;
		rom[ 23   ] = 8'h00;
		rom[ 24   ] = 8'h43;
		rom[ 25   ] = 8'h00;
		// quantization table index 0 begins
		rom[ 26   ] = 8'h10;
		rom[ 27   ] = 8'h0B;
		rom[ 28   ] = 8'h0C;
		rom[ 29   ] = 8'h0E;
		rom[ 30   ] = 8'h0C;
		rom[ 31   ] = 8'h0A;
		rom[ 32   ] = 8'h10;
		rom[ 33   ] = 8'h0E;
		rom[ 34   ] = 8'h0D;
		rom[ 35   ] = 8'h0E;
		rom[ 36   ] = 8'h12;
		rom[ 37   ] = 8'h11;
		rom[ 38   ] = 8'h10;
		rom[ 39   ] = 8'h13;
		rom[ 40   ] = 8'h18;
		rom[ 41   ] = 8'h28;
		rom[ 42   ] = 8'h1A;
		rom[ 43   ] = 8'h18;
		rom[ 44   ] = 8'h16;
		rom[ 45   ] = 8'h16;
		rom[ 46   ] = 8'h18;
		rom[ 47   ] = 8'h31;
		rom[ 48   ] = 8'h23;
		rom[ 49   ] = 8'h25;
		rom[ 50   ] = 8'h1D;
		rom[ 51   ] = 8'h28;
		rom[ 52   ] = 8'h3A;
		rom[ 53   ] = 8'h33;
		rom[ 54   ] = 8'h3D;
		rom[ 55   ] = 8'h3C;
		rom[ 56   ] = 8'h39;
		rom[ 57   ] = 8'h33;
		rom[ 58   ] = 8'h38;
		rom[ 59   ] = 8'h37;
		rom[ 60   ] = 8'h40;
		rom[ 61   ] = 8'h48;
		rom[ 62   ] = 8'h5C;
		rom[ 63   ] = 8'h4E;
		rom[ 64   ] = 8'h40;
		rom[ 65   ] = 8'h44;
		rom[ 66   ] = 8'h57;
		rom[ 67   ] = 8'h45;
		rom[ 68   ] = 8'h37;
		rom[ 69   ] = 8'h38;
		rom[ 70   ] = 8'h50;
		rom[ 71   ] = 8'h6D;
		rom[ 72   ] = 8'h51;
		rom[ 73   ] = 8'h57;
		rom[ 74   ] = 8'h5F;
		rom[ 75   ] = 8'h62;
		rom[ 76   ] = 8'h67;
		rom[ 77   ] = 8'h68;
		rom[ 78   ] = 8'h67;
		rom[ 79   ] = 8'h3E;
		rom[ 80   ] = 8'h4D;
		rom[ 81   ] = 8'h71;
		rom[ 82   ] = 8'h79;
		rom[ 83   ] = 8'h70;
		rom[ 84   ] = 8'h64;
		rom[ 85   ] = 8'h78;
		rom[ 86   ] = 8'h5C;
		rom[ 87   ] = 8'h65;
		rom[ 88   ] = 8'h67;
		rom[ 89   ] = 8'h63;
		// quantization table index 1 header begins
		rom[ 90   ] = 8'hFF;
		rom[ 91   ] = 8'hDB;
		rom[ 92   ] = 8'h00;
		rom[ 93   ] = 8'h43;
		rom[ 94   ] = 8'h01;
		// quantization table index 1 begins
		rom[ 95   ] = 8'h11;
		rom[ 96   ] = 8'h12;
		rom[ 97   ] = 8'h12;
		rom[ 98   ] = 8'h18;
		rom[ 99   ] = 8'h15;
		rom[ 100  ] = 8'h18;
		rom[ 101  ] = 8'h2F;
		rom[ 102  ] = 8'h1A;
		rom[ 103  ] = 8'h1A;
		rom[ 104  ] = 8'h2F;
		rom[ 105  ] = 8'h63;
		rom[ 106  ] = 8'h42;
		rom[ 107  ] = 8'h38;
		rom[ 108  ] = 8'h42;
		rom[ 109  ] = 8'h63;
		rom[ 110  ] = 8'h63;
		rom[ 111  ] = 8'h63;
		rom[ 112  ] = 8'h63;
		rom[ 113  ] = 8'h63;
		rom[ 114  ] = 8'h63;
		rom[ 115  ] = 8'h63;
		rom[ 116  ] = 8'h63;
		rom[ 117  ] = 8'h63;
		rom[ 118  ] = 8'h63;
		rom[ 119  ] = 8'h63;
		rom[ 120  ] = 8'h63;
		rom[ 121  ] = 8'h63;
		rom[ 122  ] = 8'h63;
		rom[ 123  ] = 8'h63;
		rom[ 124  ] = 8'h63;
		rom[ 125  ] = 8'h63;
		rom[ 126  ] = 8'h63;
		rom[ 127  ] = 8'h63;
		rom[ 128  ] = 8'h63;
		rom[ 129  ] = 8'h63;
		rom[ 130  ] = 8'h63;
		rom[ 131  ] = 8'h63;
		rom[ 132  ] = 8'h63;
		rom[ 133  ] = 8'h63;
		rom[ 134  ] = 8'h63;
		rom[ 135  ] = 8'h63;
		rom[ 136  ] = 8'h63;
		rom[ 137  ] = 8'h63;
		rom[ 138  ] = 8'h63;
		rom[ 139  ] = 8'h63;
		rom[ 140  ] = 8'h63;
		rom[ 141  ] = 8'h63;
		rom[ 142  ] = 8'h63;
		rom[ 143  ] = 8'h63;
		rom[ 144  ] = 8'h63;
		rom[ 145  ] = 8'h63;
		rom[ 146  ] = 8'h63;
		rom[ 147  ] = 8'h63;
		rom[ 148  ] = 8'h63;
		rom[ 149  ] = 8'h63;
		rom[ 150  ] = 8'h63;
		rom[ 151  ] = 8'h63;
		rom[ 152  ] = 8'h63;
		rom[ 153  ] = 8'h63;
		rom[ 154  ] = 8'h63;
		rom[ 155  ] = 8'h63;
		rom[ 156  ] = 8'h63;
		rom[ 157  ] = 8'h63;
		rom[ 158  ] = 8'h63;
		// Huffmann table header begins
		rom[ 159  ] = 8'hFF;
		rom[ 160  ] = 8'hC4;
		rom[ 161  ] = 8'h00;
		rom[ 162  ] = 8'h1F; //31-2-1 = 28
		// huffmann bits
		rom[ 163  ] = 8'h00;
		rom[ 164  ] = 8'h00;
		rom[ 165  ] = 8'h01;
		rom[ 166  ] = 8'h05;
		rom[ 167  ] = 8'h01;
		rom[ 168  ] = 8'h01;
		rom[ 169  ] = 8'h01;
		rom[ 170  ] = 8'h01;
		rom[ 171  ] = 8'h01;
		rom[ 172  ] = 8'h01;
		rom[ 173  ] = 8'h00;
		rom[ 174  ] = 8'h00;
		rom[ 175  ] = 8'h00;
		rom[ 176  ] = 8'h00;
		rom[ 177  ] = 8'h00;
		rom[ 178  ] = 8'h00;
		rom[ 179  ] = 8'h00;
		rom[ 180  ] = 8'h00;

		rom[ 181  ] = 8'h01;
		rom[ 182  ] = 8'h02;
		rom[ 183  ] = 8'h03;
		rom[ 184  ] = 8'h04;
		rom[ 185  ] = 8'h05;
		rom[ 186  ] = 8'h06;
		rom[ 187  ] = 8'h07;
		rom[ 188  ] = 8'h08;
		rom[ 189  ] = 8'h09;
		rom[ 190  ] = 8'h0A;
		rom[ 191  ] = 8'h0B;

		rom[ 192  ] = 8'hFF;
		rom[ 193  ] = 8'hC4;
		rom[ 194  ] = 8'h00;
		rom[ 195  ] = 8'h1F;
		rom[ 196  ] = 8'h01;
		rom[ 197  ] = 8'h00;
		rom[ 198  ] = 8'h03;
		rom[ 199  ] = 8'h01;
		rom[ 200  ] = 8'h01;
		rom[ 201  ] = 8'h01;
		rom[ 202  ] = 8'h01;
		rom[ 203  ] = 8'h01;
		rom[ 204  ] = 8'h01;
		rom[ 205  ] = 8'h01;
		rom[ 206  ] = 8'h01;
		rom[ 207  ] = 8'h01;
		rom[ 208  ] = 8'h00;
		rom[ 209  ] = 8'h00;
		rom[ 210  ] = 8'h00;
		rom[ 211  ] = 8'h00;
		rom[ 212  ] = 8'h00;
		rom[ 213  ] = 8'h00;
		rom[ 214  ] = 8'h01;
		rom[ 215  ] = 8'h02;
		rom[ 216  ] = 8'h03;
		rom[ 217  ] = 8'h04;
		rom[ 218  ] = 8'h05;
		rom[ 219  ] = 8'h06;
		rom[ 220  ] = 8'h07;
		rom[ 221  ] = 8'h08;
		rom[ 222  ] = 8'h09;
		rom[ 223  ] = 8'h0A;
		rom[ 224  ] = 8'h0B;

		rom[ 225  ] = 8'hFF;
		rom[ 226  ] = 8'hC4;
		rom[ 227  ] = 8'h00;
		rom[ 228  ] = 8'hB5;
		rom[ 229  ] = 8'h10;
		rom[ 230  ] = 8'h00;
		rom[ 231  ] = 8'h02;
		rom[ 232  ] = 8'h01;
		rom[ 233  ] = 8'h03;
		rom[ 234  ] = 8'h03;
		rom[ 235  ] = 8'h02;
		rom[ 236  ] = 8'h04;
		rom[ 237  ] = 8'h03;
		rom[ 238  ] = 8'h05;
		rom[ 239  ] = 8'h05;
		rom[ 240  ] = 8'h04;
		rom[ 241  ] = 8'h04;
		rom[ 242  ] = 8'h00;
		rom[ 243  ] = 8'h00;
		rom[ 244  ] = 8'h01;
		rom[ 245  ] = 8'h7D;
		rom[ 246  ] = 8'h01;
		rom[ 247  ] = 8'h02;
		rom[ 248  ] = 8'h03;
		rom[ 249  ] = 8'h00;
		rom[ 250  ] = 8'h04;
		rom[ 251  ] = 8'h11;
		rom[ 252  ] = 8'h05;
		rom[ 253  ] = 8'h12;
		rom[ 254  ] = 8'h21;
		rom[ 255  ] = 8'h31;
		rom[ 256  ] = 8'h41;
		rom[ 257  ] = 8'h06;
		rom[ 258  ] = 8'h13;
		rom[ 259  ] = 8'h51;
		rom[ 260  ] = 8'h61;
		rom[ 261  ] = 8'h07;
		rom[ 262  ] = 8'h22;
		rom[ 263  ] = 8'h71;
		rom[ 264  ] = 8'h14;
		rom[ 265  ] = 8'h32;
		rom[ 266  ] = 8'h81;
		rom[ 267  ] = 8'h91;
		rom[ 268  ] = 8'hA1;
		rom[ 269  ] = 8'h08;
		rom[ 270  ] = 8'h23;
		rom[ 271  ] = 8'h42;
		rom[ 272  ] = 8'hB1;
		rom[ 273  ] = 8'hC1;
		rom[ 274  ] = 8'h15;
		rom[ 275  ] = 8'h52;
		rom[ 276  ] = 8'hD1;
		rom[ 277  ] = 8'hF0;
		rom[ 278  ] = 8'h24;
		rom[ 279  ] = 8'h33;
		rom[ 280  ] = 8'h62;
		rom[ 281  ] = 8'h72;
		rom[ 282  ] = 8'h82;
		rom[ 283  ] = 8'h09;
		rom[ 284  ] = 8'h0A;
		rom[ 285  ] = 8'h16;
		rom[ 286  ] = 8'h17;
		rom[ 287  ] = 8'h18;
		rom[ 288  ] = 8'h19;
		rom[ 289  ] = 8'h1A;
		rom[ 290  ] = 8'h25;
		rom[ 291  ] = 8'h26;
		rom[ 292  ] = 8'h27;
		rom[ 293  ] = 8'h28;
		rom[ 294  ] = 8'h29;
		rom[ 295  ] = 8'h2A;
		rom[ 296  ] = 8'h34;
		rom[ 297  ] = 8'h35;
		rom[ 298  ] = 8'h36;
		rom[ 299  ] = 8'h37;
		rom[ 300  ] = 8'h38;
		rom[ 301  ] = 8'h39;
		rom[ 302  ] = 8'h3A;
		rom[ 303  ] = 8'h43;
		rom[ 304  ] = 8'h44;
		rom[ 305  ] = 8'h45;
		rom[ 306  ] = 8'h46;
		rom[ 307  ] = 8'h47;
		rom[ 308  ] = 8'h48;
		rom[ 309  ] = 8'h49;
		rom[ 310  ] = 8'h4A;
		rom[ 311  ] = 8'h53;
		rom[ 312  ] = 8'h54;
		rom[ 313  ] = 8'h55;
		rom[ 314  ] = 8'h56;
		rom[ 315  ] = 8'h57;
		rom[ 316  ] = 8'h58;
		rom[ 317  ] = 8'h59;
		rom[ 318  ] = 8'h5A;
		rom[ 319  ] = 8'h63;
		rom[ 320  ] = 8'h64;
		rom[ 321  ] = 8'h65;
		rom[ 322  ] = 8'h66;
		rom[ 323  ] = 8'h67;
		rom[ 324  ] = 8'h68;
		rom[ 325  ] = 8'h69;
		rom[ 326  ] = 8'h6A;
		rom[ 327  ] = 8'h73;
		rom[ 328  ] = 8'h74;
		rom[ 329  ] = 8'h75;
		rom[ 330  ] = 8'h76;
		rom[ 331  ] = 8'h77;
		rom[ 332  ] = 8'h78;
		rom[ 333  ] = 8'h79;
		rom[ 334  ] = 8'h7A;
		rom[ 335  ] = 8'h83;
		rom[ 336  ] = 8'h84;
		rom[ 337  ] = 8'h85;
		rom[ 338  ] = 8'h86;
		rom[ 339  ] = 8'h87;
		rom[ 340  ] = 8'h88;
		rom[ 341  ] = 8'h89;
		rom[ 342  ] = 8'h8A;
		rom[ 343  ] = 8'h92;
		rom[ 344  ] = 8'h93;
		rom[ 345  ] = 8'h94;
		rom[ 346  ] = 8'h95;
		rom[ 347  ] = 8'h96;
		rom[ 348  ] = 8'h97;
		rom[ 349  ] = 8'h98;
		rom[ 350  ] = 8'h99;
		rom[ 351  ] = 8'h9A;
		rom[ 352  ] = 8'hA2;
		rom[ 353  ] = 8'hA3;
		rom[ 354  ] = 8'hA4;
		rom[ 355  ] = 8'hA5;
		rom[ 356  ] = 8'hA6;
		rom[ 357  ] = 8'hA7;
		rom[ 358  ] = 8'hA8;
		rom[ 359  ] = 8'hA9;
		rom[ 360  ] = 8'hAA;
		rom[ 361  ] = 8'hB2;
		rom[ 362  ] = 8'hB3;
		rom[ 363  ] = 8'hB4;
		rom[ 364  ] = 8'hB5;
		rom[ 365  ] = 8'hB6;
		rom[ 366  ] = 8'hB7;
		rom[ 367  ] = 8'hB8;
		rom[ 368  ] = 8'hB9;
		rom[ 369  ] = 8'hBA;
		rom[ 370  ] = 8'hC2;
		rom[ 371  ] = 8'hC3;
		rom[ 372  ] = 8'hC4;
		rom[ 373  ] = 8'hC5;
		rom[ 374  ] = 8'hC6;
		rom[ 375  ] = 8'hC7;
		rom[ 376  ] = 8'hC8;
		rom[ 377  ] = 8'hC9;
		rom[ 378  ] = 8'hCA;
		rom[ 379  ] = 8'hD2;
		rom[ 380  ] = 8'hD3;
		rom[ 381  ] = 8'hD4;
		rom[ 382  ] = 8'hD5;
		rom[ 383  ] = 8'hD6;
		rom[ 384  ] = 8'hD7;
		rom[ 385  ] = 8'hD8;
		rom[ 386  ] = 8'hD9;
		rom[ 387  ] = 8'hDA;
		rom[ 388  ] = 8'hE1;
		rom[ 389  ] = 8'hE2;
		rom[ 390  ] = 8'hE3;
		rom[ 391  ] = 8'hE4;
		rom[ 392  ] = 8'hE5;
		rom[ 393  ] = 8'hE6;
		rom[ 394  ] = 8'hE7;
		rom[ 395  ] = 8'hE8;
		rom[ 396  ] = 8'hE9;
		rom[ 397  ] = 8'hEA;
		rom[ 398  ] = 8'hF1;
		rom[ 399  ] = 8'hF2;
		rom[ 400  ] = 8'hF3;
		rom[ 401  ] = 8'hF4;
		rom[ 402  ] = 8'hF5;
		rom[ 403  ] = 8'hF6;
		rom[ 404  ] = 8'hF7;
		rom[ 405  ] = 8'hF8;
		rom[ 406  ] = 8'hF9;
		rom[ 407  ] = 8'hFA;
		rom[ 408  ] = 8'hFF;
		rom[ 409  ] = 8'hC4;
		rom[ 410  ] = 8'h00;
		rom[ 411  ] = 8'hB5;
		rom[ 412  ] = 8'h11;
		rom[ 413  ] = 8'h00;
		rom[ 414  ] = 8'h02;
		rom[ 415  ] = 8'h01;
		rom[ 416  ] = 8'h02;
		rom[ 417  ] = 8'h04;
		rom[ 418  ] = 8'h04;
		rom[ 419  ] = 8'h03;
		rom[ 420  ] = 8'h04;
		rom[ 421  ] = 8'h07;
		rom[ 422  ] = 8'h05;
		rom[ 423  ] = 8'h04;
		rom[ 424  ] = 8'h04;
		rom[ 425  ] = 8'h00;
		rom[ 426  ] = 8'h01;
		rom[ 427  ] = 8'h02;
		rom[ 428  ] = 8'h77;
		rom[ 429  ] = 8'h00;
		rom[ 430  ] = 8'h01;
		rom[ 431  ] = 8'h02;
		rom[ 432  ] = 8'h03;
		rom[ 433  ] = 8'h11;
		rom[ 434  ] = 8'h04;
		rom[ 435  ] = 8'h05;
		rom[ 436  ] = 8'h21;
		rom[ 437  ] = 8'h31;
		rom[ 438  ] = 8'h06;
		rom[ 439  ] = 8'h12;
		rom[ 440  ] = 8'h41;
		rom[ 441  ] = 8'h51;
		rom[ 442  ] = 8'h07;
		rom[ 443  ] = 8'h61;
		rom[ 444  ] = 8'h71;
		rom[ 445  ] = 8'h13;
		rom[ 446  ] = 8'h22;
		rom[ 447  ] = 8'h32;
		rom[ 448  ] = 8'h81;
		rom[ 449  ] = 8'h08;
		rom[ 450  ] = 8'h14;
		rom[ 451  ] = 8'h42;
		rom[ 452  ] = 8'h91;
		rom[ 453  ] = 8'hA1;
		rom[ 454  ] = 8'hB1;
		rom[ 455  ] = 8'hC1;
		rom[ 456  ] = 8'h09;
		rom[ 457  ] = 8'h23;
		rom[ 458  ] = 8'h33;
		rom[ 459  ] = 8'h52;
		rom[ 460  ] = 8'hF0;
		rom[ 461  ] = 8'h15;
		rom[ 462  ] = 8'h62;
		rom[ 463  ] = 8'h72;
		rom[ 464  ] = 8'hD1;
		rom[ 465  ] = 8'h0A;
		rom[ 466  ] = 8'h16;
		rom[ 467  ] = 8'h24;
		rom[ 468  ] = 8'h34;
		rom[ 469  ] = 8'hE1;
		rom[ 470  ] = 8'h25;
		rom[ 471  ] = 8'hF1;
		rom[ 472  ] = 8'h17;
		rom[ 473  ] = 8'h18;
		rom[ 474  ] = 8'h19;
		rom[ 475  ] = 8'h1A;
		rom[ 476  ] = 8'h26;
		rom[ 477  ] = 8'h27;
		rom[ 478  ] = 8'h28;
		rom[ 479  ] = 8'h29;
		rom[ 480  ] = 8'h2A;
		rom[ 481  ] = 8'h35;
		rom[ 482  ] = 8'h36;
		rom[ 483  ] = 8'h37;
		rom[ 484  ] = 8'h38;
		rom[ 485  ] = 8'h39;
		rom[ 486  ] = 8'h3A;
		rom[ 487  ] = 8'h43;
		rom[ 488  ] = 8'h44;
		rom[ 489  ] = 8'h45;
		rom[ 490  ] = 8'h46;
		rom[ 491  ] = 8'h47;
		rom[ 492  ] = 8'h48;
		rom[ 493  ] = 8'h49;
		rom[ 494  ] = 8'h4A;
		rom[ 495  ] = 8'h53;
		rom[ 496  ] = 8'h54;
		rom[ 497  ] = 8'h55;
		rom[ 498  ] = 8'h56;
		rom[ 499  ] = 8'h57;
		rom[ 500  ] = 8'h58;
		rom[ 501  ] = 8'h59;
		rom[ 502  ] = 8'h5A;
		rom[ 503  ] = 8'h63;
		rom[ 504  ] = 8'h64;
		rom[ 505  ] = 8'h65;
		rom[ 506  ] = 8'h66;
		rom[ 507  ] = 8'h67;
		rom[ 508  ] = 8'h68;
		rom[ 509  ] = 8'h69;
		rom[ 510  ] = 8'h6A;
		rom[ 511  ] = 8'h73;
		rom[ 512  ] = 8'h74;
		rom[ 513  ] = 8'h75;
		rom[ 514  ] = 8'h76;
		rom[ 515  ] = 8'h77;
		rom[ 516  ] = 8'h78;
		rom[ 517  ] = 8'h79;
		rom[ 518  ] = 8'h7A;
		rom[ 519  ] = 8'h82;
		rom[ 520  ] = 8'h83;
		rom[ 521  ] = 8'h84;
		rom[ 522  ] = 8'h85;
		rom[ 523  ] = 8'h86;
		rom[ 524  ] = 8'h87;
		rom[ 525  ] = 8'h88;
		rom[ 526  ] = 8'h89;
		rom[ 527  ] = 8'h8A;
		rom[ 528  ] = 8'h92;
		rom[ 529  ] = 8'h93;
		rom[ 530  ] = 8'h94;
		rom[ 531  ] = 8'h95;
		rom[ 532  ] = 8'h96;
		rom[ 533  ] = 8'h97;
		rom[ 534  ] = 8'h98;
		rom[ 535  ] = 8'h99;
		rom[ 536  ] = 8'h9A;
		rom[ 537  ] = 8'hA2;
		rom[ 538  ] = 8'hA3;
		rom[ 539  ] = 8'hA4;
		rom[ 540  ] = 8'hA5;
		rom[ 541  ] = 8'hA6;
		rom[ 542  ] = 8'hA7;
		rom[ 543  ] = 8'hA8;
		rom[ 544  ] = 8'hA9;
		rom[ 545  ] = 8'hAA;
		rom[ 546  ] = 8'hB2;
		rom[ 547  ] = 8'hB3;
		rom[ 548  ] = 8'hB4;
		rom[ 549  ] = 8'hB5;
		rom[ 550  ] = 8'hB6;
		rom[ 551  ] = 8'hB7;
		rom[ 552  ] = 8'hB8;
		rom[ 553  ] = 8'hB9;
		rom[ 554  ] = 8'hBA;
		rom[ 555  ] = 8'hC2;
		rom[ 556  ] = 8'hC3;
		rom[ 557  ] = 8'hC4;
		rom[ 558  ] = 8'hC5;
		rom[ 559  ] = 8'hC6;
		rom[ 560  ] = 8'hC7;
		rom[ 561  ] = 8'hC8;
		rom[ 562  ] = 8'hC9;
		rom[ 563  ] = 8'hCA;
		rom[ 564  ] = 8'hD2;
		rom[ 565  ] = 8'hD3;
		rom[ 566  ] = 8'hD4;
		rom[ 567  ] = 8'hD5;
		rom[ 568  ] = 8'hD6;
		rom[ 569  ] = 8'hD7;
		rom[ 570  ] = 8'hD8;
		rom[ 571  ] = 8'hD9;
		rom[ 572  ] = 8'hDA;
		rom[ 573  ] = 8'hE2;
		rom[ 574  ] = 8'hE3;
		rom[ 575  ] = 8'hE4;
		rom[ 576  ] = 8'hE5;
		rom[ 577  ] = 8'hE6;
		rom[ 578  ] = 8'hE7;
		rom[ 579  ] = 8'hE8;
		rom[ 580  ] = 8'hE9;
		rom[ 581  ] = 8'hEA;
		rom[ 582  ] = 8'hF2;
		rom[ 583  ] = 8'hF3;
		rom[ 584  ] = 8'hF4;
		rom[ 585  ] = 8'hF5;
		rom[ 586  ] = 8'hF6;
		rom[ 587  ] = 8'hF7;
		rom[ 588  ] = 8'hF8;
		rom[ 589  ] = 8'hF9;
		rom[ 590  ] = 8'hFA;
		rom[ 591  ] = 8'hFF;
		rom[ 592  ] = 8'hDA;
		rom[ 593  ] = 8'h00;
		rom[ 594  ] = 8'h0C;
		rom[ 595  ] = 8'h03;
		rom[ 596  ] = 8'h01;
		rom[ 597  ] = 8'h00;
		rom[ 598  ] = 8'h02;
		rom[ 599  ] = 8'h11;
		rom[ 600  ] = 8'h03;
		rom[ 601  ] = 8'h11;
		rom[ 602  ] = 8'h00;
		rom[ 603  ] = 8'h3F;
		rom[ 604  ] = 8'h00;
	end
endmodule


module rom_header_qf09(
	input 				clk,
	input		[9:0]	addr,
	output reg	[7:0]	q
	);
	
	reg					[7:0]	rom [1023:0];
	always @(posedge clk) q <= rom[addr];
	initial begin
		rom[ 0    ] = 8'hFF;
		rom[ 1    ] = 8'hD8;
		rom[ 2    ] = 8'hFF;
		rom[ 3    ] = 8'hC0;
		rom[ 4    ] = 8'h00;
		rom[ 5    ] = 8'h11;
		rom[ 6    ] = 8'h08;
		rom[ 7    ] = 8'h01;
		rom[ 8    ] = 8'h20;
		rom[ 9    ] = 8'h01;
		rom[ 10   ] = 8'h60;
		rom[ 11   ] = 8'h03;
		rom[ 12   ] = 8'h01;
`ifdef YUV444_ONLY
		rom[ 13   ] = 8'h11;
`elsif YUV422_ONLY
		rom[ 13   ] = 8'h21;
`endif
		rom[ 14   ] = 8'h00;
		rom[ 15   ] = 8'h02;
		rom[ 16   ] = 8'h11;
		rom[ 17   ] = 8'h01;
		rom[ 18   ] = 8'h03;
		rom[ 19   ] = 8'h11;
		rom[ 20   ] = 8'h01;
		// quantization table index 0 header begins
		rom[ 21   ] = 8'hFF;
		rom[ 22   ] = 8'hDB;
		rom[ 23   ] = 8'h00;
		rom[ 24   ] = 8'h43;
		rom[ 25   ] = 8'h00;
		// quantization table index 0 begins
		rom[ 26   ] = 8'h03;
		rom[ 27   ] = 8'h02;
		rom[ 28   ] = 8'h02;
		rom[ 29   ] = 8'h02;
		rom[ 30   ] = 8'h02;
		rom[ 31   ] = 8'h03;
		rom[ 32   ] = 8'h03;
		rom[ 33   ] = 8'h03;
		rom[ 34   ] = 8'h03;
		rom[ 35   ] = 8'h03;
		rom[ 36   ] = 8'h05;
		rom[ 37   ] = 8'h04;
		rom[ 38   ] = 8'h03;
		rom[ 39   ] = 8'h03;
		rom[ 40   ] = 8'h04;
		rom[ 41   ] = 8'h05;
		rom[ 42   ] = 8'h04;
		rom[ 43   ] = 8'h04;
		rom[ 44   ] = 8'h05;
		rom[ 45   ] = 8'h05;
		rom[ 46   ] = 8'h08;
		rom[ 47   ] = 8'h0a;
		rom[ 48   ] = 8'h0c;
		rom[ 49   ] = 8'h08;
		rom[ 50   ] = 8'h06;
		rom[ 51   ] = 8'h07;
		rom[ 52   ] = 8'h07;
		rom[ 53   ] = 8'h0a;
		rom[ 54   ] = 8'h0e;
		rom[ 55   ] = 8'h0d;
		rom[ 56   ] = 8'h0b;
		rom[ 57   ] = 8'h0b;
		rom[ 58   ] = 8'h0a;
		rom[ 59   ] = 8'h0b;
		rom[ 60   ] = 8'h0c;
		rom[ 61   ] = 8'h0c;
		rom[ 62   ] = 8'h0b;
		rom[ 63   ] = 8'h0e;
		rom[ 64   ] = 8'h11;
		rom[ 65   ] = 8'h0e;
		rom[ 66   ] = 8'h0d;
		rom[ 67   ] = 8'h10;
		rom[ 68   ] = 8'h12;
		rom[ 69   ] = 8'h13;
		rom[ 70   ] = 8'h11;
		rom[ 71   ] = 8'h10;
		rom[ 72   ] = 8'h16;
		rom[ 73   ] = 8'h10;
		rom[ 74   ] = 8'h0b;
		rom[ 75   ] = 8'h0c;
		rom[ 76   ] = 8'h15;
		rom[ 77   ] = 8'h15;
		rom[ 78   ] = 8'h15;
		rom[ 79   ] = 8'h14;
		rom[ 80   ] = 8'h16;
		rom[ 81   ] = 8'h18;
		rom[ 82   ] = 8'h17;
		rom[ 83   ] = 8'h0f;
		rom[ 84   ] = 8'h12;
		rom[ 85   ] = 8'h18;
		rom[ 86   ] = 8'h14;
		rom[ 87   ] = 8'h15;
		rom[ 88   ] = 8'h14;
		rom[ 89   ] = 8'h14;
		// quantization table index 1 header begins
		rom[ 90   ] = 8'hFF;
		rom[ 91   ] = 8'hDB;
		rom[ 92   ] = 8'h00;
		rom[ 93   ] = 8'h43;
		rom[ 94   ] = 8'h01;
		// quantization table index 1 begins
		rom[ 95   ] = 8'h03;
		rom[ 96   ] = 8'h04;
		rom[ 97   ] = 8'h04;
		rom[ 98   ] = 8'h05;
		rom[ 99   ] = 8'h04;
		rom[ 100   ] = 8'h05;
		rom[ 101   ] = 8'h09;
		rom[ 102   ] = 8'h05;
		rom[ 103   ] = 8'h05;
		rom[ 104   ] = 8'h09;
		rom[ 105   ] = 8'h14;
		rom[ 106   ] = 8'h0d;
		rom[ 107   ] = 8'h0b;
		rom[ 108   ] = 8'h0d;
		rom[ 109   ] = 8'h14;
		rom[ 110   ] = 8'h14;
		rom[ 111   ] = 8'h14;
		rom[ 112   ] = 8'h14;
		rom[ 113   ] = 8'h14;
		rom[ 114   ] = 8'h14;
		rom[ 115   ] = 8'h14;
		rom[ 116   ] = 8'h14;
		rom[ 117   ] = 8'h14;
		rom[ 118   ] = 8'h14;
		rom[ 119   ] = 8'h14;
		rom[ 120   ] = 8'h14;
		rom[ 121   ] = 8'h14;
		rom[ 122   ] = 8'h14;
		rom[ 123   ] = 8'h14;
		rom[ 124   ] = 8'h14;
		rom[ 125   ] = 8'h14;
		rom[ 126   ] = 8'h14;
		rom[ 127   ] = 8'h14;
		rom[ 128   ] = 8'h14;
		rom[ 129   ] = 8'h14;
		rom[ 130   ] = 8'h14;
		rom[ 131   ] = 8'h14;
		rom[ 132   ] = 8'h14;
		rom[ 133   ] = 8'h14;
		rom[ 134   ] = 8'h14;
		rom[ 135   ] = 8'h14;
		rom[ 136   ] = 8'h14;
		rom[ 137   ] = 8'h14;
		rom[ 138   ] = 8'h14;
		rom[ 139   ] = 8'h14;
		rom[ 140   ] = 8'h14;
		rom[ 141   ] = 8'h14;
		rom[ 142   ] = 8'h14;
		rom[ 143   ] = 8'h14;
		rom[ 144   ] = 8'h14;
		rom[ 145   ] = 8'h14;
		rom[ 146   ] = 8'h14;
		rom[ 147   ] = 8'h14;
		rom[ 148   ] = 8'h14;
		rom[ 149   ] = 8'h14;
		rom[ 150   ] = 8'h14;
		rom[ 151   ] = 8'h14;
		rom[ 152   ] = 8'h14;
		rom[ 153   ] = 8'h14;
		rom[ 154   ] = 8'h14;
		rom[ 155   ] = 8'h14;
		rom[ 156   ] = 8'h14;
		rom[ 157   ] = 8'h14;
		rom[ 158   ] = 8'h14;
		// Huffmann table header begins
		rom[ 159  ] = 8'hFF;
		rom[ 160  ] = 8'hC4;
		rom[ 161  ] = 8'h00;
		rom[ 162  ] = 8'h1F; //31-2-1 = 28
		// huffmann bits
		rom[ 163  ] = 8'h00;
		rom[ 164  ] = 8'h00;
		rom[ 165  ] = 8'h01;
		rom[ 166  ] = 8'h05;
		rom[ 167  ] = 8'h01;
		rom[ 168  ] = 8'h01;
		rom[ 169  ] = 8'h01;
		rom[ 170  ] = 8'h01;
		rom[ 171  ] = 8'h01;
		rom[ 172  ] = 8'h01;
		rom[ 173  ] = 8'h00;
		rom[ 174  ] = 8'h00;
		rom[ 175  ] = 8'h00;
		rom[ 176  ] = 8'h00;
		rom[ 177  ] = 8'h00;
		rom[ 178  ] = 8'h00;
		rom[ 179  ] = 8'h00;
		rom[ 180  ] = 8'h00;

		rom[ 181  ] = 8'h01;
		rom[ 182  ] = 8'h02;
		rom[ 183  ] = 8'h03;
		rom[ 184  ] = 8'h04;
		rom[ 185  ] = 8'h05;
		rom[ 186  ] = 8'h06;
		rom[ 187  ] = 8'h07;
		rom[ 188  ] = 8'h08;
		rom[ 189  ] = 8'h09;
		rom[ 190  ] = 8'h0A;
		rom[ 191  ] = 8'h0B;

		rom[ 192  ] = 8'hFF;
		rom[ 193  ] = 8'hC4;
		rom[ 194  ] = 8'h00;
		rom[ 195  ] = 8'h1F;
		rom[ 196  ] = 8'h01;
		rom[ 197  ] = 8'h00;
		rom[ 198  ] = 8'h03;
		rom[ 199  ] = 8'h01;
		rom[ 200  ] = 8'h01;
		rom[ 201  ] = 8'h01;
		rom[ 202  ] = 8'h01;
		rom[ 203  ] = 8'h01;
		rom[ 204  ] = 8'h01;
		rom[ 205  ] = 8'h01;
		rom[ 206  ] = 8'h01;
		rom[ 207  ] = 8'h01;
		rom[ 208  ] = 8'h00;
		rom[ 209  ] = 8'h00;
		rom[ 210  ] = 8'h00;
		rom[ 211  ] = 8'h00;
		rom[ 212  ] = 8'h00;
		rom[ 213  ] = 8'h00;
		rom[ 214  ] = 8'h01;
		rom[ 215  ] = 8'h02;
		rom[ 216  ] = 8'h03;
		rom[ 217  ] = 8'h04;
		rom[ 218  ] = 8'h05;
		rom[ 219  ] = 8'h06;
		rom[ 220  ] = 8'h07;
		rom[ 221  ] = 8'h08;
		rom[ 222  ] = 8'h09;
		rom[ 223  ] = 8'h0A;
		rom[ 224  ] = 8'h0B;

		rom[ 225  ] = 8'hFF;
		rom[ 226  ] = 8'hC4;
		rom[ 227  ] = 8'h00;
		rom[ 228  ] = 8'hB5;
		rom[ 229  ] = 8'h10;
		rom[ 230  ] = 8'h00;
		rom[ 231  ] = 8'h02;
		rom[ 232  ] = 8'h01;
		rom[ 233  ] = 8'h03;
		rom[ 234  ] = 8'h03;
		rom[ 235  ] = 8'h02;
		rom[ 236  ] = 8'h04;
		rom[ 237  ] = 8'h03;
		rom[ 238  ] = 8'h05;
		rom[ 239  ] = 8'h05;
		rom[ 240  ] = 8'h04;
		rom[ 241  ] = 8'h04;
		rom[ 242  ] = 8'h00;
		rom[ 243  ] = 8'h00;
		rom[ 244  ] = 8'h01;
		rom[ 245  ] = 8'h7D;
		rom[ 246  ] = 8'h01;
		rom[ 247  ] = 8'h02;
		rom[ 248  ] = 8'h03;
		rom[ 249  ] = 8'h00;
		rom[ 250  ] = 8'h04;
		rom[ 251  ] = 8'h11;
		rom[ 252  ] = 8'h05;
		rom[ 253  ] = 8'h12;
		rom[ 254  ] = 8'h21;
		rom[ 255  ] = 8'h31;
		rom[ 256  ] = 8'h41;
		rom[ 257  ] = 8'h06;
		rom[ 258  ] = 8'h13;
		rom[ 259  ] = 8'h51;
		rom[ 260  ] = 8'h61;
		rom[ 261  ] = 8'h07;
		rom[ 262  ] = 8'h22;
		rom[ 263  ] = 8'h71;
		rom[ 264  ] = 8'h14;
		rom[ 265  ] = 8'h32;
		rom[ 266  ] = 8'h81;
		rom[ 267  ] = 8'h91;
		rom[ 268  ] = 8'hA1;
		rom[ 269  ] = 8'h08;
		rom[ 270  ] = 8'h23;
		rom[ 271  ] = 8'h42;
		rom[ 272  ] = 8'hB1;
		rom[ 273  ] = 8'hC1;
		rom[ 274  ] = 8'h15;
		rom[ 275  ] = 8'h52;
		rom[ 276  ] = 8'hD1;
		rom[ 277  ] = 8'hF0;
		rom[ 278  ] = 8'h24;
		rom[ 279  ] = 8'h33;
		rom[ 280  ] = 8'h62;
		rom[ 281  ] = 8'h72;
		rom[ 282  ] = 8'h82;
		rom[ 283  ] = 8'h09;
		rom[ 284  ] = 8'h0A;
		rom[ 285  ] = 8'h16;
		rom[ 286  ] = 8'h17;
		rom[ 287  ] = 8'h18;
		rom[ 288  ] = 8'h19;
		rom[ 289  ] = 8'h1A;
		rom[ 290  ] = 8'h25;
		rom[ 291  ] = 8'h26;
		rom[ 292  ] = 8'h27;
		rom[ 293  ] = 8'h28;
		rom[ 294  ] = 8'h29;
		rom[ 295  ] = 8'h2A;
		rom[ 296  ] = 8'h34;
		rom[ 297  ] = 8'h35;
		rom[ 298  ] = 8'h36;
		rom[ 299  ] = 8'h37;
		rom[ 300  ] = 8'h38;
		rom[ 301  ] = 8'h39;
		rom[ 302  ] = 8'h3A;
		rom[ 303  ] = 8'h43;
		rom[ 304  ] = 8'h44;
		rom[ 305  ] = 8'h45;
		rom[ 306  ] = 8'h46;
		rom[ 307  ] = 8'h47;
		rom[ 308  ] = 8'h48;
		rom[ 309  ] = 8'h49;
		rom[ 310  ] = 8'h4A;
		rom[ 311  ] = 8'h53;
		rom[ 312  ] = 8'h54;
		rom[ 313  ] = 8'h55;
		rom[ 314  ] = 8'h56;
		rom[ 315  ] = 8'h57;
		rom[ 316  ] = 8'h58;
		rom[ 317  ] = 8'h59;
		rom[ 318  ] = 8'h5A;
		rom[ 319  ] = 8'h63;
		rom[ 320  ] = 8'h64;
		rom[ 321  ] = 8'h65;
		rom[ 322  ] = 8'h66;
		rom[ 323  ] = 8'h67;
		rom[ 324  ] = 8'h68;
		rom[ 325  ] = 8'h69;
		rom[ 326  ] = 8'h6A;
		rom[ 327  ] = 8'h73;
		rom[ 328  ] = 8'h74;
		rom[ 329  ] = 8'h75;
		rom[ 330  ] = 8'h76;
		rom[ 331  ] = 8'h77;
		rom[ 332  ] = 8'h78;
		rom[ 333  ] = 8'h79;
		rom[ 334  ] = 8'h7A;
		rom[ 335  ] = 8'h83;
		rom[ 336  ] = 8'h84;
		rom[ 337  ] = 8'h85;
		rom[ 338  ] = 8'h86;
		rom[ 339  ] = 8'h87;
		rom[ 340  ] = 8'h88;
		rom[ 341  ] = 8'h89;
		rom[ 342  ] = 8'h8A;
		rom[ 343  ] = 8'h92;
		rom[ 344  ] = 8'h93;
		rom[ 345  ] = 8'h94;
		rom[ 346  ] = 8'h95;
		rom[ 347  ] = 8'h96;
		rom[ 348  ] = 8'h97;
		rom[ 349  ] = 8'h98;
		rom[ 350  ] = 8'h99;
		rom[ 351  ] = 8'h9A;
		rom[ 352  ] = 8'hA2;
		rom[ 353  ] = 8'hA3;
		rom[ 354  ] = 8'hA4;
		rom[ 355  ] = 8'hA5;
		rom[ 356  ] = 8'hA6;
		rom[ 357  ] = 8'hA7;
		rom[ 358  ] = 8'hA8;
		rom[ 359  ] = 8'hA9;
		rom[ 360  ] = 8'hAA;
		rom[ 361  ] = 8'hB2;
		rom[ 362  ] = 8'hB3;
		rom[ 363  ] = 8'hB4;
		rom[ 364  ] = 8'hB5;
		rom[ 365  ] = 8'hB6;
		rom[ 366  ] = 8'hB7;
		rom[ 367  ] = 8'hB8;
		rom[ 368  ] = 8'hB9;
		rom[ 369  ] = 8'hBA;
		rom[ 370  ] = 8'hC2;
		rom[ 371  ] = 8'hC3;
		rom[ 372  ] = 8'hC4;
		rom[ 373  ] = 8'hC5;
		rom[ 374  ] = 8'hC6;
		rom[ 375  ] = 8'hC7;
		rom[ 376  ] = 8'hC8;
		rom[ 377  ] = 8'hC9;
		rom[ 378  ] = 8'hCA;
		rom[ 379  ] = 8'hD2;
		rom[ 380  ] = 8'hD3;
		rom[ 381  ] = 8'hD4;
		rom[ 382  ] = 8'hD5;
		rom[ 383  ] = 8'hD6;
		rom[ 384  ] = 8'hD7;
		rom[ 385  ] = 8'hD8;
		rom[ 386  ] = 8'hD9;
		rom[ 387  ] = 8'hDA;
		rom[ 388  ] = 8'hE1;
		rom[ 389  ] = 8'hE2;
		rom[ 390  ] = 8'hE3;
		rom[ 391  ] = 8'hE4;
		rom[ 392  ] = 8'hE5;
		rom[ 393  ] = 8'hE6;
		rom[ 394  ] = 8'hE7;
		rom[ 395  ] = 8'hE8;
		rom[ 396  ] = 8'hE9;
		rom[ 397  ] = 8'hEA;
		rom[ 398  ] = 8'hF1;
		rom[ 399  ] = 8'hF2;
		rom[ 400  ] = 8'hF3;
		rom[ 401  ] = 8'hF4;
		rom[ 402  ] = 8'hF5;
		rom[ 403  ] = 8'hF6;
		rom[ 404  ] = 8'hF7;
		rom[ 405  ] = 8'hF8;
		rom[ 406  ] = 8'hF9;
		rom[ 407  ] = 8'hFA;
		rom[ 408  ] = 8'hFF;
		rom[ 409  ] = 8'hC4;
		rom[ 410  ] = 8'h00;
		rom[ 411  ] = 8'hB5;
		rom[ 412  ] = 8'h11;
		rom[ 413  ] = 8'h00;
		rom[ 414  ] = 8'h02;
		rom[ 415  ] = 8'h01;
		rom[ 416  ] = 8'h02;
		rom[ 417  ] = 8'h04;
		rom[ 418  ] = 8'h04;
		rom[ 419  ] = 8'h03;
		rom[ 420  ] = 8'h04;
		rom[ 421  ] = 8'h07;
		rom[ 422  ] = 8'h05;
		rom[ 423  ] = 8'h04;
		rom[ 424  ] = 8'h04;
		rom[ 425  ] = 8'h00;
		rom[ 426  ] = 8'h01;
		rom[ 427  ] = 8'h02;
		rom[ 428  ] = 8'h77;
		rom[ 429  ] = 8'h00;
		rom[ 430  ] = 8'h01;
		rom[ 431  ] = 8'h02;
		rom[ 432  ] = 8'h03;
		rom[ 433  ] = 8'h11;
		rom[ 434  ] = 8'h04;
		rom[ 435  ] = 8'h05;
		rom[ 436  ] = 8'h21;
		rom[ 437  ] = 8'h31;
		rom[ 438  ] = 8'h06;
		rom[ 439  ] = 8'h12;
		rom[ 440  ] = 8'h41;
		rom[ 441  ] = 8'h51;
		rom[ 442  ] = 8'h07;
		rom[ 443  ] = 8'h61;
		rom[ 444  ] = 8'h71;
		rom[ 445  ] = 8'h13;
		rom[ 446  ] = 8'h22;
		rom[ 447  ] = 8'h32;
		rom[ 448  ] = 8'h81;
		rom[ 449  ] = 8'h08;
		rom[ 450  ] = 8'h14;
		rom[ 451  ] = 8'h42;
		rom[ 452  ] = 8'h91;
		rom[ 453  ] = 8'hA1;
		rom[ 454  ] = 8'hB1;
		rom[ 455  ] = 8'hC1;
		rom[ 456  ] = 8'h09;
		rom[ 457  ] = 8'h23;
		rom[ 458  ] = 8'h33;
		rom[ 459  ] = 8'h52;
		rom[ 460  ] = 8'hF0;
		rom[ 461  ] = 8'h15;
		rom[ 462  ] = 8'h62;
		rom[ 463  ] = 8'h72;
		rom[ 464  ] = 8'hD1;
		rom[ 465  ] = 8'h0A;
		rom[ 466  ] = 8'h16;
		rom[ 467  ] = 8'h24;
		rom[ 468  ] = 8'h34;
		rom[ 469  ] = 8'hE1;
		rom[ 470  ] = 8'h25;
		rom[ 471  ] = 8'hF1;
		rom[ 472  ] = 8'h17;
		rom[ 473  ] = 8'h18;
		rom[ 474  ] = 8'h19;
		rom[ 475  ] = 8'h1A;
		rom[ 476  ] = 8'h26;
		rom[ 477  ] = 8'h27;
		rom[ 478  ] = 8'h28;
		rom[ 479  ] = 8'h29;
		rom[ 480  ] = 8'h2A;
		rom[ 481  ] = 8'h35;
		rom[ 482  ] = 8'h36;
		rom[ 483  ] = 8'h37;
		rom[ 484  ] = 8'h38;
		rom[ 485  ] = 8'h39;
		rom[ 486  ] = 8'h3A;
		rom[ 487  ] = 8'h43;
		rom[ 488  ] = 8'h44;
		rom[ 489  ] = 8'h45;
		rom[ 490  ] = 8'h46;
		rom[ 491  ] = 8'h47;
		rom[ 492  ] = 8'h48;
		rom[ 493  ] = 8'h49;
		rom[ 494  ] = 8'h4A;
		rom[ 495  ] = 8'h53;
		rom[ 496  ] = 8'h54;
		rom[ 497  ] = 8'h55;
		rom[ 498  ] = 8'h56;
		rom[ 499  ] = 8'h57;
		rom[ 500  ] = 8'h58;
		rom[ 501  ] = 8'h59;
		rom[ 502  ] = 8'h5A;
		rom[ 503  ] = 8'h63;
		rom[ 504  ] = 8'h64;
		rom[ 505  ] = 8'h65;
		rom[ 506  ] = 8'h66;
		rom[ 507  ] = 8'h67;
		rom[ 508  ] = 8'h68;
		rom[ 509  ] = 8'h69;
		rom[ 510  ] = 8'h6A;
		rom[ 511  ] = 8'h73;
		rom[ 512  ] = 8'h74;
		rom[ 513  ] = 8'h75;
		rom[ 514  ] = 8'h76;
		rom[ 515  ] = 8'h77;
		rom[ 516  ] = 8'h78;
		rom[ 517  ] = 8'h79;
		rom[ 518  ] = 8'h7A;
		rom[ 519  ] = 8'h82;
		rom[ 520  ] = 8'h83;
		rom[ 521  ] = 8'h84;
		rom[ 522  ] = 8'h85;
		rom[ 523  ] = 8'h86;
		rom[ 524  ] = 8'h87;
		rom[ 525  ] = 8'h88;
		rom[ 526  ] = 8'h89;
		rom[ 527  ] = 8'h8A;
		rom[ 528  ] = 8'h92;
		rom[ 529  ] = 8'h93;
		rom[ 530  ] = 8'h94;
		rom[ 531  ] = 8'h95;
		rom[ 532  ] = 8'h96;
		rom[ 533  ] = 8'h97;
		rom[ 534  ] = 8'h98;
		rom[ 535  ] = 8'h99;
		rom[ 536  ] = 8'h9A;
		rom[ 537  ] = 8'hA2;
		rom[ 538  ] = 8'hA3;
		rom[ 539  ] = 8'hA4;
		rom[ 540  ] = 8'hA5;
		rom[ 541  ] = 8'hA6;
		rom[ 542  ] = 8'hA7;
		rom[ 543  ] = 8'hA8;
		rom[ 544  ] = 8'hA9;
		rom[ 545  ] = 8'hAA;
		rom[ 546  ] = 8'hB2;
		rom[ 547  ] = 8'hB3;
		rom[ 548  ] = 8'hB4;
		rom[ 549  ] = 8'hB5;
		rom[ 550  ] = 8'hB6;
		rom[ 551  ] = 8'hB7;
		rom[ 552  ] = 8'hB8;
		rom[ 553  ] = 8'hB9;
		rom[ 554  ] = 8'hBA;
		rom[ 555  ] = 8'hC2;
		rom[ 556  ] = 8'hC3;
		rom[ 557  ] = 8'hC4;
		rom[ 558  ] = 8'hC5;
		rom[ 559  ] = 8'hC6;
		rom[ 560  ] = 8'hC7;
		rom[ 561  ] = 8'hC8;
		rom[ 562  ] = 8'hC9;
		rom[ 563  ] = 8'hCA;
		rom[ 564  ] = 8'hD2;
		rom[ 565  ] = 8'hD3;
		rom[ 566  ] = 8'hD4;
		rom[ 567  ] = 8'hD5;
		rom[ 568  ] = 8'hD6;
		rom[ 569  ] = 8'hD7;
		rom[ 570  ] = 8'hD8;
		rom[ 571  ] = 8'hD9;
		rom[ 572  ] = 8'hDA;
		rom[ 573  ] = 8'hE2;
		rom[ 574  ] = 8'hE3;
		rom[ 575  ] = 8'hE4;
		rom[ 576  ] = 8'hE5;
		rom[ 577  ] = 8'hE6;
		rom[ 578  ] = 8'hE7;
		rom[ 579  ] = 8'hE8;
		rom[ 580  ] = 8'hE9;
		rom[ 581  ] = 8'hEA;
		rom[ 582  ] = 8'hF2;
		rom[ 583  ] = 8'hF3;
		rom[ 584  ] = 8'hF4;
		rom[ 585  ] = 8'hF5;
		rom[ 586  ] = 8'hF6;
		rom[ 587  ] = 8'hF7;
		rom[ 588  ] = 8'hF8;
		rom[ 589  ] = 8'hF9;
		rom[ 590  ] = 8'hFA;
		rom[ 591  ] = 8'hFF;
		rom[ 592  ] = 8'hDA;
		rom[ 593  ] = 8'h00;
		rom[ 594  ] = 8'h0C;
		rom[ 595  ] = 8'h03;
		rom[ 596  ] = 8'h01;
		rom[ 597  ] = 8'h00;
		rom[ 598  ] = 8'h02;
		rom[ 599  ] = 8'h11;
		rom[ 600  ] = 8'h03;
		rom[ 601  ] = 8'h11;
		rom[ 602  ] = 8'h00;
		rom[ 603  ] = 8'h3F;
		rom[ 604  ] = 8'h00;
	end
endmodule